module vdummy

pub fn zero() int {
	return 0
}
